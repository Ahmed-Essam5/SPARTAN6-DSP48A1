module DSP48A1_Project (a,b,d,c,carryin,m,p,carryout,carryoutf,clk,opmode,cea,ceb,cec,cecarryin,ced,cem,ceopmode,cep,rsta,rstb,rstc,rstcarryin,rstd,rstm,rstopmode,rstp,bcin,bcout,pcin,pcout);

/*PARAMETERS*/
	parameter A0REG=0;
	parameter A1REG=1;
	parameter B0REG=0;
	parameter B1REG=1;
	parameter CREG=1;
	parameter DREG=1;
	parameter MREG=1;
	parameter PREG=1;
	parameter CARRYINREG=1;
	parameter CARRYOUTREG=1;
	parameter OPMODEREG=1;

	parameter CARRYINSEL="OPMODE5"; //select bet. CARRYIN or OPMODE5 or tie
	parameter B_INPUT="DIRECT"; //DIRECT(B) ,CASCADE(BCIN), tie
	parameter RSTTYPE="SYNC"; //SYNC, ASYNC

/*INPUT PORTS*/
/*DATA*/
	input [17:0]a,b,d;
	input [47:0]c;
	input carryin;
	output [35:0]m;
	output [47:0]p;
	output carryout,carryoutf;

/*CONTROL*/
	input clk;
	input [7:0]opmode;

/*ENABLE*/
	input cea,ceb,cec,cecarryin,ced,cem,ceopmode,cep; //cecarryin for carry in/out

/*RESET*/
	input rsta,rstb,rstc,rstcarryin,rstd,rstm,rstopmode,rstp; //same in rstcarryin

/*CASCADE*/
	input [17:0]bcin;
	output [17:0]bcout;
	input [47:0]pcin;
	output [47:0]pcout;

//WIRES
	wire [17:0]wa0,wa1,wb0,wb1,wd;
	wire [47:0]wc;
	wire wcarryin;
	wire [7:0]wopmode;
	wire [17:0] Pre_Adder_Subtractor;
	wire [47:0] Post_Adder_Subtractor;
	wire wcarryout_prev;
	wire [35:0] wm;
	wire [17:0] b00;
	wire carryin00;

	wire [35:0] wm00;
	assign wm00=(wa1 * wb1);

//SELECTIONS
	reg [47:0] X,Z;

//INSTATIATION
	//DSP48A1_Project_reg #(.WIDTH(), .REGISTER(), .RSTTYPE()) dut (clk,enable,rst,in,out);
	DSP48A1_Project_reg #(.WIDTH(18), .REGISTER(A0REG), .RSTTYPE(RSTTYPE)) duta0 (clk,cea,rsta,a,wa0);
	DSP48A1_Project_reg #(.WIDTH(18), .REGISTER(A1REG), .RSTTYPE(RSTTYPE)) duta1 (clk,cea,rsta,wa0,wa1);
	DSP48A1_Project_reg #(.WIDTH(18), .REGISTER(B0REG), .RSTTYPE(RSTTYPE)) dutb0 (clk,ceb,rstb,b00,wb0);
	DSP48A1_Project_reg #(.WIDTH(18), .REGISTER(B1REG), .RSTTYPE(RSTTYPE)) dutb1 (clk,ceb,rstb,((wopmode[4])?Pre_Adder_Subtractor:wb0),wb1);
	DSP48A1_Project_reg #(.WIDTH(18), .REGISTER(DREG), .RSTTYPE(RSTTYPE)) dutd (clk,ced,rstd,d,wd);
	DSP48A1_Project_reg #(.WIDTH(48), .REGISTER(CREG), .RSTTYPE(RSTTYPE)) dutc (clk,cec,rstc,c,wc);
	DSP48A1_Project_reg #(.WIDTH(1), .REGISTER(CARRYINREG), .RSTTYPE(RSTTYPE)) dutcarryin (clk,cecarryin,rstcarryin,carryin00,wcarryin);
	DSP48A1_Project_reg #(.WIDTH(36), .REGISTER(MREG), .RSTTYPE(RSTTYPE)) dutm (clk,cem,rstm,wm00,wm);
	DSP48A1_Project_reg #(.WIDTH(8), .REGISTER(OPMODEREG), .RSTTYPE(RSTTYPE)) dutopmode (clk,ceopmode,rstopmode,opmode,wopmode);
	DSP48A1_Project_reg #(.WIDTH(48), .REGISTER(PREG), .RSTTYPE(RSTTYPE)) dutP (clk,cep,rstp,Post_Adder_Subtractor,p);
	DSP48A1_Project_reg #(.WIDTH(1), .REGISTER(CARRYOUTREG), .RSTTYPE(RSTTYPE)) dutacarryout (clk,cecarryin,rstcarryin,wcarryout_prev,carryout);

	assign b00=(B_INPUT=="DIRECT")? b:(B_INPUT=="CASCADE")? bcin: 0;
	assign carryin00=(CARRYINSEL=="OPMODE5")? wopmode[5]:(CARRYINSEL=="CARRYIN")? carryin: 0;
//Pre_Adder_Subtractor
	assign Pre_Adder_Subtractor=(wopmode[6])?(wd - wb0):(wd + wb0);
//Post_Adder_Subtractor
	assign {wcarryout_prev,Post_Adder_Subtractor}=(wopmode[7])?(Z - (X + wcarryin)):(Z + X + wcarryin);
	assign carryoutf=carryout;
	assign pcout=p;
	assign bcout=wb1;
//m_buffer
	genvar i;
	generate
		for (i = 0;i <36;i=i+1) begin
			buf (m[i],wm[i]);
		end
	endgenerate

//X
	always @(*) begin
		case (wopmode[1:0])
			2'b00:X=0;
			2'b01:X=wm;
			2'b10:X=p;
			2'b11:X={d[11:0],a[17:0],b[17:0]};
		endcase
	end
//Z
	always @(*) begin
		case (wopmode[3:2])
			2'b00:Z=0;
			2'b01:Z=pcin;
			2'b10:Z=p;
			2'b11:Z=wc;
		endcase
	end

endmodule